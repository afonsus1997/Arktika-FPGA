module top (
    input CLK,
    output D13
    );
  
  assign D13 = 1;

endmodule
